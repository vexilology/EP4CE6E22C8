module signal((* chip_pin = "58" *)input X,
              (* chip_pin = "72" *)output Y);

  assign Y = X;

endmodule
